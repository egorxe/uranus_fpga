library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;
    use ieee.std_logic_unsigned.all;
    use ieee.std_logic_textio.all;

use STD.textio.all;

library fpgalib;
    use fpgalib.fpga_pkg.all;

package fpga_tb_pkg is

--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
--                                  CONSTANTS
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------

constant CFG_CLK_PERIOD     : time := 1000 ns;

--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
--                                  TYPES
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------


--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
--                                  FUNCTIONS
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------

end fpga_tb_pkg;

package body fpga_tb_pkg is

end fpga_tb_pkg;
