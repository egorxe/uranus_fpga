module fpga_memory (
    input        clk_i,
     
    input        ce_a_i,
    input  [6:0] addr_a_i,
    output [7:0] data_a_o,
    
    input        we_b_i,
    input  [6:0] addr_b_i,
    input  [7:0] data_b_i
);

// blackbox

endmodule